library verilog;
use verilog.vl_types.all;
entity cnt10_38_vlg_vec_tst is
end cnt10_38_vlg_vec_tst;
