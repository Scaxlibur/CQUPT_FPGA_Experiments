library verilog;
use verilog.vl_types.all;
entity m100_38_vlg_check_tst is
    port(
        clkout38        : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end m100_38_vlg_check_tst;
