library verilog;
use verilog.vl_types.all;
entity mux3_38_vlg_check_tst is
    port(
        bell38          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end mux3_38_vlg_check_tst;
