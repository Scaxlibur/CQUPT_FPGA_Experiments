library verilog;
use verilog.vl_types.all;
entity m100_38 is
    port(
        clkout38        : out    vl_logic;
        clk38           : in     vl_logic
    );
end m100_38;
