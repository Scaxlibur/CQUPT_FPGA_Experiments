library verilog;
use verilog.vl_types.all;
entity \123\ is
    port(
        q               : out    vl_logic_vector(3 downto 0);
        clk             : in     vl_logic
    );
end \123\;
