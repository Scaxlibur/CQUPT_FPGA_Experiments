library verilog;
use verilog.vl_types.all;
entity m100_38_vlg_sample_tst is
    port(
        clk38           : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end m100_38_vlg_sample_tst;
