library verilog;
use verilog.vl_types.all;
entity cnt10_38 is
    port(
        q38             : out    vl_logic_vector(2 downto 0);
        CLK_IN38        : in     vl_logic
    );
end cnt10_38;
