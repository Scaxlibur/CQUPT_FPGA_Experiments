library verilog;
use verilog.vl_types.all;
entity cnt10_38_vlg_sample_tst is
    port(
        CLK_IN38        : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end cnt10_38_vlg_sample_tst;
